module AHB2APB_BNridge(


) ;



endmodule